// DE2_115_SOPC.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module DE2_115_SOPC (
		output wire        altpll_sys,                   //            c0_out_clk.clk
		output wire        altpll_io,                    //            c2_out_clk.clk
		input  wire        clk_50,                       //         clk_50_clk_in.clk
		input  wire        reset_n,                      //   clk_50_clk_in_reset.reset_n
		output wire [31:0] mouse_data_EXPORT_DATA,       //            mouse_data.EXPORT_DATA
		output wire        altpll_sdram,                 //                pll_c1.clk
		output wire        altpll_25,                    //                pll_c3.clk
		output wire        locked_from_the_pll,          //    pll_locked_conduit.export
		output wire        phasedone_from_the_pll,       // pll_phasedone_conduit.export
		output wire [12:0] zs_addr_from_the_sdram,       //            sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,         //                      .ba
		output wire        zs_cas_n_from_the_sdram,      //                      .cas_n
		output wire        zs_cke_from_the_sdram,        //                      .cke
		output wire        zs_cs_n_from_the_sdram,       //                      .cs_n
		inout  wire [31:0] zs_dq_to_and_from_the_sdram,  //                      .dq
		output wire [3:0]  zs_dqm_from_the_sdram,        //                      .dqm
		output wire        zs_ras_n_from_the_sdram,      //                      .ras_n
		output wire        zs_we_n_from_the_sdram,       //                      .we_n
		inout  wire [15:0] SRAM_DQ_to_and_from_the_sram, //      sram_conduit_end.DQ
		output wire [19:0] SRAM_ADDR_from_the_sram,      //                      .ADDR
		output wire        SRAM_UB_n_from_the_sram,      //                      .UB_n
		output wire        SRAM_LB_n_from_the_sram,      //                      .LB_n
		output wire        SRAM_WE_n_from_the_sram,      //                      .WE_n
		output wire        SRAM_CE_n_from_the_sram,      //                      .CE_n
		output wire        SRAM_OE_n_from_the_sram,      //                      .OE_n
		inout  wire [15:0] usb_conduit_end_DATA,         //       usb_conduit_end.DATA
		output wire [1:0]  usb_conduit_end_ADDR,         //                      .ADDR
		output wire        usb_conduit_end_RD_N,         //                      .RD_N
		output wire        usb_conduit_end_WR_N,         //                      .WR_N
		output wire        usb_conduit_end_CS_N,         //                      .CS_N
		output wire        usb_conduit_end_RST_N,        //                      .RST_N
		input  wire        usb_conduit_end_INT           //                      .INT
	);

	wire  [31:0] cpu_data_master_readdata;                                     // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                  // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                  // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                      // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                   // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                         // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                        // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                    // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                              // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                           // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                               // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                  // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                         // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_mouse_core_remake_0_mouse_slave_chipselect; // mm_interconnect_0:mouse_core_remake_0_MOUSE_SLAVE_chipselect -> mouse_core_remake_0:AVL_CS
	wire  [31:0] mm_interconnect_0_mouse_core_remake_0_mouse_slave_readdata;   // mouse_core_remake_0:AVL_READDATA -> mm_interconnect_0:mouse_core_remake_0_MOUSE_SLAVE_readdata
	wire   [3:0] mm_interconnect_0_mouse_core_remake_0_mouse_slave_address;    // mm_interconnect_0:mouse_core_remake_0_MOUSE_SLAVE_address -> mouse_core_remake_0:AVL_ADDR
	wire         mm_interconnect_0_mouse_core_remake_0_mouse_slave_read;       // mm_interconnect_0:mouse_core_remake_0_MOUSE_SLAVE_read -> mouse_core_remake_0:AVL_READ
	wire   [3:0] mm_interconnect_0_mouse_core_remake_0_mouse_slave_byteenable; // mm_interconnect_0:mouse_core_remake_0_MOUSE_SLAVE_byteenable -> mouse_core_remake_0:AVL_BYTE_EN
	wire         mm_interconnect_0_mouse_core_remake_0_mouse_slave_write;      // mm_interconnect_0:mouse_core_remake_0_MOUSE_SLAVE_write -> mouse_core_remake_0:AVL_WRITE
	wire  [31:0] mm_interconnect_0_mouse_core_remake_0_mouse_slave_writedata;  // mm_interconnect_0:mouse_core_remake_0_MOUSE_SLAVE_writedata -> mouse_core_remake_0:AVL_WRITEDATA
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_sram_avalon_slave_chipselect;               // mm_interconnect_0:sram_avalon_slave_chipselect -> sram:s_chipselect_n
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_readdata;                 // sram:s_readdata -> mm_interconnect_0:sram_avalon_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_slave_address;                  // mm_interconnect_0:sram_avalon_slave_address -> sram:s_address
	wire         mm_interconnect_0_sram_avalon_slave_read;                     // mm_interconnect_0:sram_avalon_slave_read -> sram:s_read_n
	wire   [1:0] mm_interconnect_0_sram_avalon_slave_byteenable;               // mm_interconnect_0:sram_avalon_slave_byteenable -> sram:s_byteenable_n
	wire         mm_interconnect_0_sram_avalon_slave_write;                    // mm_interconnect_0:sram_avalon_slave_write -> sram:s_write_n
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_writedata;                // mm_interconnect_0:sram_avalon_slave_writedata -> sram:s_writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;             // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;          // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;          // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;              // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                 // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;           // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;            // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                     // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                      // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                         // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                        // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                    // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;              // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;           // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;           // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire  [21:0] mm_interconnect_0_clock_crossing_io_s0_address;               // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                  // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;            // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;         // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                 // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;             // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;            // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                        // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                          // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                       // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                           // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                              // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                        // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                     // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                             // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                         // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_stamp_s1_chipselect;                  // mm_interconnect_0:timer_stamp_s1_chipselect -> timer_stamp:chipselect
	wire  [15:0] mm_interconnect_0_timer_stamp_s1_readdata;                    // timer_stamp:readdata -> mm_interconnect_0:timer_stamp_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_stamp_s1_address;                     // mm_interconnect_0:timer_stamp_s1_address -> timer_stamp:address
	wire         mm_interconnect_0_timer_stamp_s1_write;                       // mm_interconnect_0:timer_stamp_s1_write -> timer_stamp:write_n
	wire  [15:0] mm_interconnect_0_timer_stamp_s1_writedata;                   // mm_interconnect_0:timer_stamp_s1_writedata -> timer_stamp:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                        // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                          // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                           // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                             // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                         // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         clock_crossing_io_m0_waitrequest;                             // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [31:0] clock_crossing_io_m0_readdata;                                // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                             // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire  [21:0] clock_crossing_io_m0_address;                                 // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire         clock_crossing_io_m0_read;                                    // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire   [3:0] clock_crossing_io_m0_byteenable;                              // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                           // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [31:0] clock_crossing_io_m0_writedata;                               // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                   // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire   [0:0] clock_crossing_io_m0_burstcount;                              // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;               // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_cy7c67200_if_0_hpi_chipselect;              // mm_interconnect_1:CY7C67200_IF_0_hpi_chipselect -> CY7C67200_IF_0:iCS_N
	wire  [31:0] mm_interconnect_1_cy7c67200_if_0_hpi_readdata;                // CY7C67200_IF_0:oDATA -> mm_interconnect_1:CY7C67200_IF_0_hpi_readdata
	wire   [1:0] mm_interconnect_1_cy7c67200_if_0_hpi_address;                 // mm_interconnect_1:CY7C67200_IF_0_hpi_address -> CY7C67200_IF_0:iADDR
	wire         mm_interconnect_1_cy7c67200_if_0_hpi_read;                    // mm_interconnect_1:CY7C67200_IF_0_hpi_read -> CY7C67200_IF_0:iRD_N
	wire         mm_interconnect_1_cy7c67200_if_0_hpi_write;                   // mm_interconnect_1:CY7C67200_IF_0_hpi_write -> CY7C67200_IF_0:iWR_N
	wire  [31:0] mm_interconnect_1_cy7c67200_if_0_hpi_writedata;               // mm_interconnect_1:CY7C67200_IF_0_hpi_writedata -> CY7C67200_IF_0:iDATA
	wire         irq_mapper_receiver2_irq;                                     // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                     // timer_stamp:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_d_irq_irq;                                                // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_receiver0_irq;                                     // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                // CY7C67200_IF_0:oINT -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                     // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                            // timer:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [CY7C67200_IF_0:iRST_N, clock_crossing_io:m0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_0:timer_reset_reset_bridge_in_reset_reset, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, sysid:reset_n, timer:reset_n]
	wire         cpu_jtag_debug_module_reset_reset;                            // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [clock_crossing_io:s0_reset, cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sram:reset_n, timer_stamp:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, mouse_core_remake_0:RESET, pll:reset]

	CY7C67200_IF cy7c67200_if_0 (
		.oDATA     (mm_interconnect_1_cy7c67200_if_0_hpi_readdata),    //              hpi.readdata
		.iADDR     (mm_interconnect_1_cy7c67200_if_0_hpi_address),     //                 .address
		.iRD_N     (~mm_interconnect_1_cy7c67200_if_0_hpi_read),       //                 .read_n
		.iWR_N     (~mm_interconnect_1_cy7c67200_if_0_hpi_write),      //                 .write_n
		.iCS_N     (~mm_interconnect_1_cy7c67200_if_0_hpi_chipselect), //                 .chipselect_n
		.iDATA     (mm_interconnect_1_cy7c67200_if_0_hpi_writedata),   //                 .writedata
		.iCLK      (altpll_io),                                        //       clock_sink.clk
		.iRST_N    (~rst_controller_reset_out_reset),                  // clock_sink_reset.reset_n
		.oINT      (irq_synchronizer_receiver_irq),                    // interrupt_sender.irq
		.HPI_DATA  (usb_conduit_end_DATA),                             //      conduit_end.export
		.HPI_ADDR  (usb_conduit_end_ADDR),                             //                 .export
		.HPI_RD_N  (usb_conduit_end_RD_N),                             //                 .export
		.HPI_WR_N  (usb_conduit_end_WR_N),                             //                 .export
		.HPI_CS_N  (usb_conduit_end_CS_N),                             //                 .export
		.HPI_RST_N (usb_conduit_end_RST_N),                            //                 .export
		.HPI_INT   (usb_conduit_end_INT)                               //                 .export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (22),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_io),                                            //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (altpll_sys),                                           //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_SOPC_cpu cpu (
		.clk                                   (altpll_sys),                                          //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE2_115_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_sys),                                                //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	avalon_mouse_interface mouse_core_remake_0 (
		.AVL_ADDR      (mm_interconnect_0_mouse_core_remake_0_mouse_slave_address),    // MOUSE_SLAVE.address
		.AVL_CS        (mm_interconnect_0_mouse_core_remake_0_mouse_slave_chipselect), //            .chipselect
		.AVL_BYTE_EN   (mm_interconnect_0_mouse_core_remake_0_mouse_slave_byteenable), //            .byteenable
		.AVL_READ      (mm_interconnect_0_mouse_core_remake_0_mouse_slave_read),       //            .read
		.AVL_READDATA  (mm_interconnect_0_mouse_core_remake_0_mouse_slave_readdata),   //            .readdata
		.AVL_WRITE     (mm_interconnect_0_mouse_core_remake_0_mouse_slave_write),      //            .write
		.AVL_WRITEDATA (mm_interconnect_0_mouse_core_remake_0_mouse_slave_writedata),  //            .writedata
		.EXPORT_DATA   (mouse_data_EXPORT_DATA),                                       // EXPORT_DATA.EXPORT_DATA
		.CLK           (clk_50),                                                       //         CLK.clk
		.RESET         (rst_controller_002_reset_out_reset)                            //       RESET.reset
	);

	DE2_115_SOPC_pll pll (
		.clk       (clk_50),                                    //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (altpll_sys),                                //                    c0.clk
		.c1        (altpll_sdram),                              //                    c1.clk
		.c2        (altpll_io),                                 //                    c2.clk
		.c3        (altpll_25),                                 //                    c3.clk
		.locked    (locked_from_the_pll),                       //        locked_conduit.export
		.phasedone (phasedone_from_the_pll)                     //     phasedone_conduit.export
	);

	DE2_115_SOPC_sdram sdram (
		.clk            (altpll_sys),                               //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	TERASIC_SRAM #(
		.DATA_BITS (16),
		.ADDR_BITS (20)
	) sram (
		.clk            (altpll_sys),                                      //       clock_reset.clk
		.reset_n        (~rst_controller_001_reset_out_reset),             // clock_reset_reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_sram_avalon_slave_chipselect), //      avalon_slave.chipselect_n
		.s_write_n      (~mm_interconnect_0_sram_avalon_slave_write),      //                  .write_n
		.s_address      (mm_interconnect_0_sram_avalon_slave_address),     //                  .address
		.s_read_n       (~mm_interconnect_0_sram_avalon_slave_read),       //                  .read_n
		.s_writedata    (mm_interconnect_0_sram_avalon_slave_writedata),   //                  .writedata
		.s_readdata     (mm_interconnect_0_sram_avalon_slave_readdata),    //                  .readdata
		.s_byteenable_n (~mm_interconnect_0_sram_avalon_slave_byteenable), //                  .byteenable_n
		.SRAM_DQ        (SRAM_DQ_to_and_from_the_sram),                    //       conduit_end.export
		.SRAM_ADDR      (SRAM_ADDR_from_the_sram),                         //                  .export
		.SRAM_UB_n      (SRAM_UB_n_from_the_sram),                         //                  .export
		.SRAM_LB_n      (SRAM_LB_n_from_the_sram),                         //                  .export
		.SRAM_WE_n      (SRAM_WE_n_from_the_sram),                         //                  .export
		.SRAM_CE_n      (SRAM_CE_n_from_the_sram),                         //                  .export
		.SRAM_OE_n      (SRAM_OE_n_from_the_sram)                          //                  .export
	);

	DE2_115_SOPC_sysid sysid (
		.clock    (altpll_io),                                      //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE2_115_SOPC_timer timer (
		.clk        (altpll_io),                             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)      //   irq.irq
	);

	DE2_115_SOPC_timer_stamp timer_stamp (
		.clk        (altpll_sys),                                  //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_stamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_stamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_stamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_stamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_stamp_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                     //   irq.irq
	);

	DE2_115_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                        (clk_50),                                                       //                                      clk_50_clk.clk
		.pll_c0_clk                                            (altpll_sys),                                                   //                                          pll_c0.clk
		.pll_c2_clk                                            (altpll_io),                                                    //                                          pll_c2.clk
		.cpu_reset_n_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                           //               cpu_reset_n_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                           // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.timer_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                               //               timer_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                      //                                 cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                                  //                                                .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                                   //                                                .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                         //                                                .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                                     //                                                .readdata
		.cpu_data_master_readdatavalid                         (cpu_data_master_readdatavalid),                                //                                                .readdatavalid
		.cpu_data_master_write                                 (cpu_data_master_write),                                        //                                                .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                                    //                                                .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                                  //                                                .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                               //                          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                           //                                                .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                                  //                                                .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                              //                                                .readdata
		.cpu_instruction_master_readdatavalid                  (cpu_instruction_master_readdatavalid),                         //                                                .readdatavalid
		.clock_crossing_io_s0_address                          (mm_interconnect_0_clock_crossing_io_s0_address),               //                            clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                            (mm_interconnect_0_clock_crossing_io_s0_write),                 //                                                .write
		.clock_crossing_io_s0_read                             (mm_interconnect_0_clock_crossing_io_s0_read),                  //                                                .read
		.clock_crossing_io_s0_readdata                         (mm_interconnect_0_clock_crossing_io_s0_readdata),              //                                                .readdata
		.clock_crossing_io_s0_writedata                        (mm_interconnect_0_clock_crossing_io_s0_writedata),             //                                                .writedata
		.clock_crossing_io_s0_burstcount                       (mm_interconnect_0_clock_crossing_io_s0_burstcount),            //                                                .burstcount
		.clock_crossing_io_s0_byteenable                       (mm_interconnect_0_clock_crossing_io_s0_byteenable),            //                                                .byteenable
		.clock_crossing_io_s0_readdatavalid                    (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),         //                                                .readdatavalid
		.clock_crossing_io_s0_waitrequest                      (mm_interconnect_0_clock_crossing_io_s0_waitrequest),           //                                                .waitrequest
		.clock_crossing_io_s0_debugaccess                      (mm_interconnect_0_clock_crossing_io_s0_debugaccess),           //                                                .debugaccess
		.cpu_jtag_debug_module_address                         (mm_interconnect_0_cpu_jtag_debug_module_address),              //                           cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                           (mm_interconnect_0_cpu_jtag_debug_module_write),                //                                                .write
		.cpu_jtag_debug_module_read                            (mm_interconnect_0_cpu_jtag_debug_module_read),                 //                                                .read
		.cpu_jtag_debug_module_readdata                        (mm_interconnect_0_cpu_jtag_debug_module_readdata),             //                                                .readdata
		.cpu_jtag_debug_module_writedata                       (mm_interconnect_0_cpu_jtag_debug_module_writedata),            //                                                .writedata
		.cpu_jtag_debug_module_byteenable                      (mm_interconnect_0_cpu_jtag_debug_module_byteenable),           //                                                .byteenable
		.cpu_jtag_debug_module_waitrequest                     (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),          //                                                .waitrequest
		.cpu_jtag_debug_module_debugaccess                     (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),          //                                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                                .chipselect
		.mouse_core_remake_0_MOUSE_SLAVE_address               (mm_interconnect_0_mouse_core_remake_0_mouse_slave_address),    //                 mouse_core_remake_0_MOUSE_SLAVE.address
		.mouse_core_remake_0_MOUSE_SLAVE_write                 (mm_interconnect_0_mouse_core_remake_0_mouse_slave_write),      //                                                .write
		.mouse_core_remake_0_MOUSE_SLAVE_read                  (mm_interconnect_0_mouse_core_remake_0_mouse_slave_read),       //                                                .read
		.mouse_core_remake_0_MOUSE_SLAVE_readdata              (mm_interconnect_0_mouse_core_remake_0_mouse_slave_readdata),   //                                                .readdata
		.mouse_core_remake_0_MOUSE_SLAVE_writedata             (mm_interconnect_0_mouse_core_remake_0_mouse_slave_writedata),  //                                                .writedata
		.mouse_core_remake_0_MOUSE_SLAVE_byteenable            (mm_interconnect_0_mouse_core_remake_0_mouse_slave_byteenable), //                                                .byteenable
		.mouse_core_remake_0_MOUSE_SLAVE_chipselect            (mm_interconnect_0_mouse_core_remake_0_mouse_slave_chipselect), //                                                .chipselect
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                      //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                        //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                         //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                     //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                    //                                                .writedata
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                           //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                             //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                              //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                          //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                         //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                        //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                     //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                       //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect),                        //                                                .chipselect
		.sram_avalon_slave_address                             (mm_interconnect_0_sram_avalon_slave_address),                  //                               sram_avalon_slave.address
		.sram_avalon_slave_write                               (mm_interconnect_0_sram_avalon_slave_write),                    //                                                .write
		.sram_avalon_slave_read                                (mm_interconnect_0_sram_avalon_slave_read),                     //                                                .read
		.sram_avalon_slave_readdata                            (mm_interconnect_0_sram_avalon_slave_readdata),                 //                                                .readdata
		.sram_avalon_slave_writedata                           (mm_interconnect_0_sram_avalon_slave_writedata),                //                                                .writedata
		.sram_avalon_slave_byteenable                          (mm_interconnect_0_sram_avalon_slave_byteenable),               //                                                .byteenable
		.sram_avalon_slave_chipselect                          (mm_interconnect_0_sram_avalon_slave_chipselect),               //                                                .chipselect
		.timer_s1_address                                      (mm_interconnect_0_timer_s1_address),                           //                                        timer_s1.address
		.timer_s1_write                                        (mm_interconnect_0_timer_s1_write),                             //                                                .write
		.timer_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                          //                                                .readdata
		.timer_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                         //                                                .writedata
		.timer_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect),                        //                                                .chipselect
		.timer_stamp_s1_address                                (mm_interconnect_0_timer_stamp_s1_address),                     //                                  timer_stamp_s1.address
		.timer_stamp_s1_write                                  (mm_interconnect_0_timer_stamp_s1_write),                       //                                                .write
		.timer_stamp_s1_readdata                               (mm_interconnect_0_timer_stamp_s1_readdata),                    //                                                .readdata
		.timer_stamp_s1_writedata                              (mm_interconnect_0_timer_stamp_s1_writedata),                   //                                                .writedata
		.timer_stamp_s1_chipselect                             (mm_interconnect_0_timer_stamp_s1_chipselect)                   //                                                .chipselect
	);

	DE2_115_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.pll_c2_clk                                             (altpll_io),                                       //                                           pll_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                  // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                    //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),                //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                 //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                 //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                       //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                   //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),              //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                      //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                  //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),                //                                                 .debugaccess
		.CY7C67200_IF_0_hpi_address                             (mm_interconnect_1_cy7c67200_if_0_hpi_address),    //                               CY7C67200_IF_0_hpi.address
		.CY7C67200_IF_0_hpi_write                               (mm_interconnect_1_cy7c67200_if_0_hpi_write),      //                                                 .write
		.CY7C67200_IF_0_hpi_read                                (mm_interconnect_1_cy7c67200_if_0_hpi_read),       //                                                 .read
		.CY7C67200_IF_0_hpi_readdata                            (mm_interconnect_1_cy7c67200_if_0_hpi_readdata),   //                                                 .readdata
		.CY7C67200_IF_0_hpi_writedata                           (mm_interconnect_1_cy7c67200_if_0_hpi_writedata),  //                                                 .writedata
		.CY7C67200_IF_0_hpi_chipselect                          (mm_interconnect_1_cy7c67200_if_0_hpi_chipselect), //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),   //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata)   //                                                 .readdata
	);

	DE2_115_SOPC_irq_mapper irq_mapper (
		.clk           (altpll_sys),                         //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                          // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (altpll_io),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (altpll_sys),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
